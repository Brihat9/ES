LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY mux2to1 IS PORT (
	SEL, I1, I2: IN STD_LOGIC;
	O: OUT STD_LOGIC
);
END mux2to1;

ARCHITECTURE dataflow OF mux2to1 IS
BEGIN
	WITH (NOT SEL AND I1) OR (SEL AND I2) SELECT
		O <= 	'1' WHEN '1',
				'0' WHEN '0',
				'0' WHEN OTHERS;
END dataflow;